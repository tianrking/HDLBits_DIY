//https://hdlbits.01xz.net/wiki/Wire

module top_module( input in, output out );
    assign out = in;
endmodule
